:))))))))
